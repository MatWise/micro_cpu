entity micro_cpu_tb is
end entity micro_cpu_tb;
