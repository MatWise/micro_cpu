entity micro_cpu_synth is
end entity micro_cpu_synth;
